LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

ENTITY decoder4_16 IS
	PORT(	    x	           :	IN		STD_LOGIC_VECTOR(3 DOWNTO 0);
	          ena          :   IN		STD_LOGIC;
			    y	           :	OUT 	STD_LOGIC_VECTOR(15 DOWNTO 0));
END ENTITY decoder4_16;
-------------------------------------------------------------
ARCHITECTURE functional OF decoder4_16 IS

SIGNAL x1 : STD_LOGIC_VECTOR(4 DOWNTO 0);

BEGIN
	
	x1 <= ena & x;
	
	y <= "0000000000000001" WHEN (x1 = "10000") ELSE 
	     "0000000000000010" WHEN (x1 = "10001") ELSE
		  "0000000000000100" WHEN (x1 = "10010") ELSE
		  "0000000000001000" WHEN (x1 = "10011") ELSE
		  "0000000000010000" WHEN (x1 = "10100") ELSE
		  "0000000000100000" WHEN (x1 = "10101") ELSE
		  "0000000001000000" WHEN (x1 = "10110") ELSE
		  "0000000010000000" WHEN (x1 = "10111") ELSE 
		  "0000000100000000" WHEN (x1 = "11000") ELSE 
	     "0000001000000000" WHEN (x1 = "11001") ELSE
		  "0000010000000000" WHEN (x1 = "11010") ELSE
		  "0000100000000000" WHEN (x1 = "11011") ELSE
		  "0001000000000000" WHEN (x1 = "11100") ELSE
		  "0010000000000000" WHEN (x1 = "11101") ELSE
		  "0100000000000000" WHEN (x1 = "11110") ELSE
		  "1000000000000000" WHEN (x1 = "11111") ELSE
		  "0000000000000000";
				  
END ARCHITECTURE functional;