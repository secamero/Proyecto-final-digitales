LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
--------------------------------------------------------------
ENTITY print_in_matrix_tb IS
END ENTITY print_in_matrix_tb;
---------------------------------------------------------------
ARCHITECTURE testbench OF print_in_matrix_tb IS

SIGNAL  clk_tb  : STD_LOGIC := '0';
SIGNAL rst_tb : STD_LOGIC := '1';
SIGNAL position_tb : STD_LOGIC_VECTOR(127 DOWNTO 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
SIGNAL filas_tb : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
SIGNAL cols1_tb : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
SIGNAL cols2_tb : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";

BEGIN

  clk_tb <= (NOT clk_tb) AFTER 10ns;
  rst_tb <= '0' AFTER 20ns;
  
--  position_tb <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" AFTER 100ns,
--                 "10000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000" AFTER 200ns,
--					  "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001" AFTER 300ns;
  
  print : ENTITY work.print_in_matrix
  PORT MAP( clk       => clk_tb,
				rst       => rst_tb,
				position  => position_tb,
            filas_out => filas_tb,
		      cols1_out => cols1_tb,
		      cols2_out => cols2_tb);
 
END ARCHITECTURE testbench; 
