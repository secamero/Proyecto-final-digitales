--LIBRARY IEEE;
--USE IEEE.std_logic_1164.all;
--USE IEEE.numeric_std.all;
--ENTITY printing IS
--  PORT (
--   
--    ROWS_IN_1  : IN  STD_LOGIC_VECTOR(0 TO 2);
--    ROWS_OUT_1 : OUT STD_LOGIC_VECTOR(0 TO 7);
--	 
--	 COLS_IN_1  : IN  STD_LOGIC_VECTOR(0 TO 127);
--	 COLS_OUT_1 : OUT STD_LOGIC_VECTOR(0 TO 15);
--	 clk			: IN	STD_LOGIC
--  );
--END ENTITY printing;
--
--ARCHITECTURE Functional OF printing IS
--
--  SIGNAL ROWS : STD_LOGIC_VECTOR(0 TO 7);
--  SIGNAL COLS : STD_LOGIC_VECTOR(0 TO 15);
--  
--BEGIN
--			
--        Encoder: ENTITY work.Mtx_Encoder
--        PORT MAP (
--		COLS_IN_0  => COLS_IN_1(0 TO 15),
--		COLS_IN_1  => COLS_IN_1(16 TO 31),
--		COLS_IN_2  => COLS_IN_1(32 TO 47),
--		COLS_IN_3  => COLS_IN_1(48 TO 63),
--		COLS_IN_4  => COLS_IN_1(64 TO 79),
--		COLS_IN_5  => COLS_IN_1(80 TO 95),
--		COLS_IN_6  => COLS_IN_1(96 TO 111),
--		COLS_IN_7  => COLS_IN_1(112 TO 127),
--		COLS_OUT   => COLS,
--      
--		ROWS_IN => ROWS_IN_1,
--		ROWS_OUT => ROWS
--        );
--		  
--  PROCESS (clk)
--  BEGIN
--    IF clk = '1' THEN
--		ROWS_OUT_1 <= ROWS;
--		COLS_OUT_1 <= COLS;
--    END IF;
--  END PROCESS;
--END ARCHITECTURE Functional;